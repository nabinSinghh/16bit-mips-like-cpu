// Top-level 16-bit CPU
// Supports: LHI, LLI, ADD, ADDI, LD, ST, HALT
// ISA: 8 registers (R0..R7), word-addressed 16-bit memory

module cpu_top (
    input  logic clk,
    input  logic reset,
    output logic halted
);

 /* 1. registers for the PC and 2. Instruction Fetch from IMEM */
    logic [15:0] pc, pc_next;
    logic  pc_en;
    logic [15:0] instr;


 /*pc module instantiation*/
    pc u_pc (
        .clk    (clk),
        .reset  (reset),
        .en     (pc_en),
        .pc_next(pc_next),
        .pc     (pc)
    );

 /*imem module instantiation*/
    imem u_imem (
        .addr (pc),  
        .data (instr)  //the 16bit instruction fetched from imem stored in instr register at cpu_top level
    );  //so we will use this 16 bit instr for decoding of the instruction, see below

 /* 3. Registers initialized for the Instruction Decode Fields */
    logic [3:0] opcode;
    logic [2:0] rs, rt, rd, funct3;
    logic [5:0] imm6;
    logic [7:0] imm8;

 //Decode instruction registers assigned
    assign opcode = instr[15:12];  //4 MSB of the instr - opcode
    assign rs = instr[11:9];  // then the further 3 bits(11:9) - source register-1
    assign rt = instr[8:6];  //next 3 bits (8:6) - source register-2/or dest for I-type
    assign rd = instr[5:3];  //dest register for R-type
    assign funct3 = instr[2:0]; //3 LSBs for R-type functtion - function

 //Immediate registers assigned, for both I-type and LHI/LLI
    assign imm6 = instr[5:0];  //normal LSB 6-bit immediate for I-type, instr[5:0]
    assign imm8 = instr[8:1];  //for LHI/LLI instructions(8 bits from instr[8:1])

 //sign-extend 6-bit immediate
    logic [15:0] imm6_sext; //sign-extended for normal I type, for immediate ALU, or offset for LD/ST or branch address
    assign imm6_sext = {{10{imm6[5]}}, imm6};  //10 0s or 1s based on sign 6th bit[5], so, sign extended to 16 bits

    //zero-extend 6-bit immediate (for ANDI / ORI)
    //for these instructions, upper 10 bits are all 0, lower 6 bits are imm6
    logic [15:0] imm6_zext;   //[15:6] = 0, [5:0] = imm6
    assign imm6_zext = {10'b0000000000, imm6};  
        //thus, imm6_sext and imm6_zext are defined at cpu_top level, and ready to be used by the I-type instructions
    //final immediate to be used by ALU (based on control signal from control unit)

 //4. Control registers defined for the CONTROL UNIT
 //these control flags/signals/1bit registers will be assigned/generated by the control unit based on opcode and funct3
 //thus, u_control will control all the muxes, based on the opcode and funct3 of the instruction
    logic reg_write;    //to write on to any of the 7 registers(r1 to r7, r0 is always 0)
    logic mem_read;     //to read from data memory(dmem)
    logic mem_write;    //to write to data memory(dmem)
    logic mem_to_reg;   //to select data memory output for writeback
    logic alu_src_imm;  //to select immediate as ALU source

    logic is_rtype;     //flag as R-type instruction
    logic is_li_type;   //flag for LHI/LLI instruction
    logic is_lhi;       //flag for LHI instruction
    logic is_lli;       //flag for LLI instruction

    //branch type flags from control unit
    logic is_beq;
    logic is_bne;
    logic is_blt;
    logic is_bge;

    logic halt;         //#####(very importatnt)  HALT signal from control

    //J-type: CALL / RET
    logic is_call;   //CALL target
    logic is_ret;    //RET

    logic is_imm_zero_ext_flag; //1bit flag to tell whether to use zero-extended(1) or sign-extended(0) imm6 for ALU

  
  //*control unit instantiation*//
  //*this unit is very important as it will generate all the control signals based on opcode and funct3*//
    control u_control (
        .opcode     (opcode),
        .funct3     (funct3),
        .reg_write  (reg_write),
        .mem_read   (mem_read),
        .mem_write  (mem_write),
        .mem_to_reg (mem_to_reg),
        .alu_src_imm (alu_src_imm),
        .is_imm_zero_ext_flag (is_imm_zero_ext_flag),
        .is_rtype   (is_rtype),
        .is_li_type (is_li_type),
        .is_lhi     (is_lhi),
        .is_lli     (is_lli),
        .halt       (halt),

        //new branch outputs from control
        .is_beq (is_beq),
        .is_bne (is_bne),
        .is_blt (is_blt),
        .is_bge (is_bge), 

        // J-type
        .is_call (is_call),
        .is_ret  (is_ret)
    );


    //FOR THE final immediate(16 bit) that goes into ALU B input when alu_src_imm = 1
    //control unit will decide whether to use sign-extended or zero-extended form
    logic [15:0] imm6_final; //16bit immediate to be used by ALU

    //for ANDI/ORI: 1 = use zero-extended imm6, 0 = use sign-extended
    //logic is_imm_zero_ext_flag;  //1bit flag from control unit, to tell if we need zero-extended(when 1) or sign-extended imm6(when 0)

    //choose which version of imm6 to use based on control signal is_imm_zero_ext_flag
    //is_imm_zero_ext_flag = 0 -> use sign-extended (ADDI, LD, ST, branches)
    //is_imm_zero_ext_flag = 1 -> use zero-extended (ANDI, ORI)
    always_comb 
    begin
        if (is_imm_zero_ext_flag)
            imm6_final = imm6_zext;  //use zero-extended version when is_imm_zero_ext_flag = 1
        else
            imm6_final = imm6_sext;  //else use sign-extended version(i.e. is_imm_zero_ext_flag = 0)
    end



 //4. Registers (out of r0 to r7, which three goes into the regfile.sv module) is defined
 //ra1, ra2, and wa are not data/registers, but the (3bit) identifiers/addresses/indices to identify which registers to access(read/write) by regfile.sv
 // and these addresses(ra1, ra2, wa) get their value from rs, rt, rd after the instruction decode (done above by cpu_top.sv)
    logic [2:0] ra1, ra2, wa; //3-bit (for 8 registers) to identify(from r0-r7) which registers to read(rs, rt) /write(rd(R-type) or rt(I-type))
    //thus, these ra1, ra2, and wa decides which one will behave as rs, rd, rt respectively from (r0 to r7)
 //for R-type, ra1 will decide whihc to be rs, ra2 will identify which to be rt, wa will decide which to be rd for R-type
 //for I-type, 
 //for ADDI/LD, ra2 is unused by the ALU (immediate is used instead). For ST/branches, ra2 = Rt is used as the second source.
  
    logic [15:0] rd1, rd2;  //to load data[16 bit] decoded by regfile (from the addresses ra1 and ra2 respectively), ready to send to alu as input A and B
    //the above are outputs from the regfile.sv module, which gives the 16bit data stored in the registers, to be used by alu/dmem

    //but below is the input, reverse of the above rd1 and rd2, this(16bit data) is given as input to regfile.sv to write into one of the registers at wa address
    logic [15:0] wd;  //writeback data[16 bit] got from alum/dmem/li_unit to write into one of the regfile(R1-R7) at address defined by wa

 // Decide which registers to read/write based on instruction type
 //in ohter words, which addresses(3 bit) to give into the ports of regfile.sv module, as rs
    always_comb 
    begin
        // By Defaults it would be for normal I-type (ADDI, ANDI, ORI, LD, ST, branches)
        //ra1 = Rs (base/source)
        //ra2 = Rt (second source for ST / branches)
        //wa  = Rt (destination for ADDI/ANDI/ORI/LD)
        ra1 = rs; //for all I type instructions, rs is the first source, so ra1 gets rs
        ra2 = rt;  //for ST and branches, rt is the second source, in other I type cases, ra2 getting rt doesn't harm(simply unused)
        wa  = rt;  //for all I type instructions, rt is the destination, so wa gets rt

        //for ohter types of instructions, we might need different assignments
        //for e.g. R-type will have wa = rd, (not rt), 
        //LHI/LLI will have ra2 = 3'd0 (unused) and so on shown in the below
        if (is_rtype) begin
            // R-type: rd = ALU(rs, rt)
            ra1 = rs;   // ALU input A = rs
            ra2 = rt;   // ALU input B = rt
            wa  = rd;   // destination = rd
        end
else if (is_li_type) begin
    // LHI/LLI: dest = Rs (bits [11:9]), old value also from Rs
    ra1 = 3'd0;      // unused
    ra2 = rs;        // rd2 = old Rs (used as old Rt in li_unit)
    wa  = rs;        // write back into Rs
end
        else if (is_call) begin
            // CALL target:
            //  LR (R7) <- PC+1, PC <- target
            //  no useful register reads, just write LR
            ra1 = 3'd0;    // unused
            ra2 = 3'd0;    // unused
            wa  = 3'b111;  // LR = R7
        end
        else if (is_ret) begin
            // RET:
            //  PC <- LR (R7)
            //  only need to read LR; no register writes
            ra1 = 3'b111;  // read LR into rd1
            ra2 = 3'd0;    // unused
            wa  = 3'd0;    // don't care (reg_write = 0 for RET)
        end
    end


 //finally after all the definitions above, we can instantiate the regfile, alu, dmem, li_unit, and writeback mux
 /***** regfile instantiation*****/
 //this takes the 1bit input reg_write/we, 3bit ra1, ra2, wa, and gets the 16bit data outputs rd1 and rd2 for to send to alu and dmem
 //or else it takes 16bit wd input from (alu, dmem, li_unit) to write into the register file, to write at wa address
    regfile u_regfile (
        .clk (clk),
        .we  (reg_write), //input-reg_write:1bit (assigned from control unit) goes into the we(write enable) of regfile
        .ra1 (ra1),    //[input-address:3bit] read address 1, assigned from above logic (cpu_top), 
        .ra2 (ra2),  //[input-address:3bit] read address 2, assigned from above logic (cpu_top)
        .wa  (wa),  //[input-address:3bit] write address, assigned from above logic (cpu_top), could differ for R-type and I-type
        .wd  (wd),//[input-data:16bit] write data, will be assigned later after alu, dmem, li_unit instantiation
        
        .rd1 (rd1),  // [output-data:16bit] read data 1, output from regfile, goes to alu input A
        .rd2 (rd2)  // [output-data:16bit] read data 2, output from regfile, goes to alu input B or dmem write data
    );



 //5.  ALU registers defined and alu instantiation
    logic [15:0] alu_a, alu_b, alu_y;  //16 bit inputs are stored in internal registers alu_a and alu_b, output in alu_y
    logic  alu_z, alu_lt_s;
    assign alu_a = rd1;  //get from the output of regfile rd1, (normal rs/rd1)
    assign alu_b = (alu_src_imm) ? imm6_final : rd2;
    //if alu_src_imm = 1, ALU B gets immediate (sign- or zero-extended), else ALU B gets rd2 from regfile
    //if is_imm_zero_ext_flag = 1, imm6_final = zero-extended imm6, else imm6_final = sign-extended imm6

 //thus, what will be inputs(alu_a, alu_b) and output(alu_y) of alu are finalized above in the cpu_top.sv
    alu u_alu (
        .A      (alu_a),  //finalized(by default) first alu input(16bit) goes to the alu input A port
        .B      (alu_b),   //finalized second alu input(16bit - either immediate or rd2) goes to the alu input B port
        .opcode (opcode),
        .funct3 (funct3),
        .Y      (alu_y),  //output (Y port from alu) is stored in the alu_y register at the cpu_top level
        .Z      (alu_z),  //1bit zero flag output(Z port) from alu stored in alu_z register at cpu_top level
        .LT_s   (alu_lt_s) //1bit signed less-than flag output(LT_s port) from alu stored in alu_lt_s register at cpu_top level
    );

    
 //6. Data memory registers defined and dmem instantiation
    logic [15:0] mem_rdata;

    dmem u_dmem (
        .clk   (clk),
        .addr  (alu_y),  //[input:16bit] address from ALU (base + offset), stored at alu_y (at cpu_top level) goes into the addr port of dmem
        .wdata (rd2),  //[input:16bit] data from the register file(rd2) to store into dmem, goes into the wdata port of dmem
        .we    (mem_write),//[input:1bit] we/write enable signal from control unit goes into the we port of dmem
        .re    (mem_read), //[input:1bit] re/read enable signal from control unit goes into the re port of dmem
        .rdata (mem_rdata) //[output:16bit] data loaded from dmem(using mem[alu_y/addr]) goes into mem_rdata register at cpu_top level 
    );                           //this mem_rdata will be used to writeback in the regfile.sv at address wa



//the writeback data(wd) to regfile.sv is decided by a mux, which selects from alu_y, mem_rdata, or pc_plus1(for CALL), or li_value(for LHI/LLI)
 //based on the control signals is_call, is_lhi/is_lli, mem_to_reg
    //thus, we need to define li_unit first to get the li_value for LHI/LLI instructions


 //7. Branch comparison logic (for BEQ, BNE, BLT, BGE)
 //these use the values already read from the register file (rd1 = Rs, rd2 = Rt)
    logic br_eq;   //1 if Rs == Rt
    logic br_lt;   //1 if Rs < Rt (signed)
    logic take_branch;

    assign br_eq = (rd1 == rd2);
    assign br_lt = ($signed(rd1) < $signed(rd2));

 //decide whether the branch is taken based on opcode-type from control
    always_comb begin
        take_branch = 1'b0; //default branch not taken

        //only one of these is expected to be 1 for a given instruction
        if (is_beq && br_eq)  //both signals, (is_beq from control and br_eq from alu comparison) should be 1
            take_branch = 1'b1;  // as soon the condition meets, take the branch
        else if (is_bne && !br_eq)  //is_bne from control should be 1 and br_eq from alu comparison should be 0
            take_branch = 1'b1;  //takes the branch, when both rd1 and rd2 are not equal
        else if (is_blt && br_lt)  //is_blt from control should be 1 and br_lt from alu comparison should be 1
            take_branch = 1'b1;
        else if (is_bge && !br_lt)  //is_bge from control should be 1 and br_lt from alu comparison should be 0
            take_branch = 1'b1;
    end

  //8. li_unit instantiation
   // LHI / LLI value generator
    logic [15:0] li_value;

    li_unit u_li (
        .is_lhi   (is_lhi),  //1bit signal from control unit
        .is_lli   (is_lli),  //1bit signal from control unit
        .imm8     (imm8),    //[input:8bit] immediate value from instruction
        .old_rt   (rd2),      // rd2 at the cpu_top level holds Rt when is_li_type = 1
        .li_value (li_value)  //[output:16bit] generated LHI/LLI value
    );


 //9. PC Next Logic
 //PC+1 and branch target address (PC+1+sign-extended offset)
    logic [15:0] pc_plus1;
    logic [15:0] branch_target;
    logic [15:0] call_target;

    //for the nomral next pc calculation, pc = pc + 1
    assign pc_plus1     = pc + 16'd1;

    //branch target address calculation, pc = pc + 1 + imm6_sext
    assign branch_target = pc_plus1 + imm6_sext;

    // J-type target address for CALL: instr[11:0] is the absolute word address
    assign call_target = {4'b0000, instr[11:0]};  //so, 4096 word address space, can access upto 4096 different instructions


 //10. Writeback Mux
    // Writeback mux section is only for what to get into the wd(16 bit write data) to the regfile.sv module at wa address
 //here, when wd at cpu_top level gets its value from alu_y, mem_rdata, li_value, or pc_plus1 
  //based on the control signals, simultaneously, wa(write address of register) at cpu_top level is already defined above
  //thus, finally regfile.sv gets both wd and wa to write into the register file
    always_comb begin
        if (is_call) begin
            wd = pc_plus1;  //CALL: LR gets PC+1
        end else if (is_lhi || is_lli) begin
            wd = li_value;  //LHI/LLI: writeback from li_unit
        end else if (mem_to_reg) begin
            wd = mem_rdata;  //writeback from memory
        end else begin
            wd = alu_y;  //DEFAULT: wd in cpu_top gets alu_y
        end
    end



 //11. HALT / PC enable logic
    logic halted_r;

    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            halted_r <= 1'b0;
        end else if (halt) begin
            halted_r <= 1'b1;
        end
    end


    assign halted  = halted_r;
    assign pc_en   = ~halted_r;

 //12. Next PC value:
    // - CALL:     jump to absolute target
    // - RET:      jump to LR (R7)
    // - branch:   PC+1+imm6 when taken
    // - default:  PC+1
    assign pc_next = (is_call) ? call_target : (is_ret) ? rd1 : (take_branch) ? branch_target : pc_plus1; 
    // rd1 holds LR when is_ret = 1   
endmodule